// sdram.v

// Generated using ACDS version 13.1 162 at 2017.12.25.22:43:06

`timescale 1 ps / 1 ps
module sdram (
		input  wire        clk_clk,                  //             clk.clk
		input  wire        reset_reset_n,            //           reset.reset_n
		input  wire        read_sdram_read_en,       //      read_sdram.read_en
		output wire [15:0] read_sdram_data,          //                .data
		input  wire [31:0] read_sdram_addr,          //                .addr
		output wire        read_sdram_dev_idle,      //                .dev_idle
		output wire        read_sdram_data_avalid,   //                .data_avalid
		input  wire        write_sdram_2_write_en,   //   write_sdram_2.write_en
		input  wire [15:0] write_sdram_2_data,       //                .data
		input  wire [31:0] write_sdram_2_addr,       //                .addr
		output wire        write_sdram_2_dev_idle,   //                .dev_idle
		input  wire        write_sdram_2_1_write_en, // write_sdram_2_1.write_en
		input  wire [15:0] write_sdram_2_1_data,     //                .data
		input  wire [31:0] write_sdram_2_1_addr,     //                .addr
		output wire        write_sdram_2_1_dev_idle, //                .dev_idle
		input  wire        write_sdram_0_write_en,   //   write_sdram_0.write_en
		input  wire [15:0] write_sdram_0_data,       //                .data
		input  wire [31:0] write_sdram_0_addr,       //                .addr
		output wire        write_sdram_0_dev_idle,   //                .dev_idle
		output wire [11:0] sdram_wire_addr,          //      sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,            //                .ba
		output wire        sdram_wire_cas_n,         //                .cas_n
		output wire        sdram_wire_cke,           //                .cke
		output wire        sdram_wire_cs_n,          //                .cs_n
		inout  wire [15:0] sdram_wire_dq,            //                .dq
		output wire [1:0]  sdram_wire_dqm,           //                .dqm
		output wire        sdram_wire_ras_n,         //                .ras_n
		output wire        sdram_wire_we_n           //                .we_n
	);

	wire   [7:0] write_sdram_burst_0_avalon_master_burstcount;  // write_sdram_burst_0:master_burstcount -> mm_interconnect_0:write_sdram_burst_0_avalon_master_burstcount
	wire         write_sdram_burst_0_avalon_master_waitrequest; // mm_interconnect_0:write_sdram_burst_0_avalon_master_waitrequest -> write_sdram_burst_0:master_waitequest
	wire  [15:0] write_sdram_burst_0_avalon_master_writedata;   // write_sdram_burst_0:master_writedata -> mm_interconnect_0:write_sdram_burst_0_avalon_master_writedata
	wire  [31:0] write_sdram_burst_0_avalon_master_address;     // write_sdram_burst_0:master_address -> mm_interconnect_0:write_sdram_burst_0_avalon_master_address
	wire         write_sdram_burst_0_avalon_master_write;       // write_sdram_burst_0:master_write -> mm_interconnect_0:write_sdram_burst_0_avalon_master_write
	wire   [1:0] write_sdram_burst_0_avalon_master_byteenable;  // write_sdram_burst_0:master_byteenable -> mm_interconnect_0:write_sdram_burst_0_avalon_master_byteenable
	wire   [7:0] write_sdram_burst_1_avalon_master_burstcount;  // write_sdram_burst_1:master_burstcount -> mm_interconnect_0:write_sdram_burst_1_avalon_master_burstcount
	wire         write_sdram_burst_1_avalon_master_waitrequest; // mm_interconnect_0:write_sdram_burst_1_avalon_master_waitrequest -> write_sdram_burst_1:master_waitequest
	wire  [15:0] write_sdram_burst_1_avalon_master_writedata;   // write_sdram_burst_1:master_writedata -> mm_interconnect_0:write_sdram_burst_1_avalon_master_writedata
	wire  [31:0] write_sdram_burst_1_avalon_master_address;     // write_sdram_burst_1:master_address -> mm_interconnect_0:write_sdram_burst_1_avalon_master_address
	wire         write_sdram_burst_1_avalon_master_write;       // write_sdram_burst_1:master_write -> mm_interconnect_0:write_sdram_burst_1_avalon_master_write
	wire   [1:0] write_sdram_burst_1_avalon_master_byteenable;  // write_sdram_burst_1:master_byteenable -> mm_interconnect_0:write_sdram_burst_1_avalon_master_byteenable
	wire         read_sdram_0_avalon_master_waitrequest;        // mm_interconnect_0:read_sdram_0_avalon_master_waitrequest -> read_sdram_0:master_waitequest
	wire  [31:0] read_sdram_0_avalon_master_address;            // read_sdram_0:master_address -> mm_interconnect_0:read_sdram_0_avalon_master_address
	wire         read_sdram_0_avalon_master_read;               // read_sdram_0:master_read -> mm_interconnect_0:read_sdram_0_avalon_master_read
	wire  [15:0] read_sdram_0_avalon_master_readdata;           // mm_interconnect_0:read_sdram_0_avalon_master_readdata -> read_sdram_0:master_readdata
	wire   [1:0] read_sdram_0_avalon_master_byteenable;         // read_sdram_0:master_byteenable -> mm_interconnect_0:read_sdram_0_avalon_master_byteenable
	wire         read_sdram_0_avalon_master_readdatavalid;      // mm_interconnect_0:read_sdram_0_avalon_master_readdatavalid -> read_sdram_0:master_readdatavalid
	wire         mm_interconnect_0_sdram_s1_waitrequest;        // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;          // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [21:0] mm_interconnect_0_sdram_s1_address;            // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;         // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;              // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;               // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;           // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;      // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;         // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire   [7:0] write_sdram_burst_2_avalon_master_burstcount;  // write_sdram_burst_2:master_burstcount -> mm_interconnect_0:write_sdram_burst_2_avalon_master_burstcount
	wire         write_sdram_burst_2_avalon_master_waitrequest; // mm_interconnect_0:write_sdram_burst_2_avalon_master_waitrequest -> write_sdram_burst_2:master_waitequest
	wire  [15:0] write_sdram_burst_2_avalon_master_writedata;   // write_sdram_burst_2:master_writedata -> mm_interconnect_0:write_sdram_burst_2_avalon_master_writedata
	wire  [31:0] write_sdram_burst_2_avalon_master_address;     // write_sdram_burst_2:master_address -> mm_interconnect_0:write_sdram_burst_2_avalon_master_address
	wire         write_sdram_burst_2_avalon_master_write;       // write_sdram_burst_2:master_write -> mm_interconnect_0:write_sdram_burst_2_avalon_master_write
	wire   [1:0] write_sdram_burst_2_avalon_master_byteenable;  // write_sdram_burst_2:master_byteenable -> mm_interconnect_0:write_sdram_burst_2_avalon_master_byteenable
	wire         rst_controller_reset_out_reset;                // rst_controller:reset_out -> [mm_interconnect_0:read_sdram_0_reset_reset_bridge_in_reset_reset, read_sdram_0:reset_n, sdram:reset_n, write_sdram_burst_0:reset_n, write_sdram_burst_1:reset_n, write_sdram_burst_2:reset_n]

	sdram_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	READ_SDRAM #(
		.IDLE    (4'b0000),
		.START   (4'b0001),
		.READING (4'b0010),
		.FINISH  (4'b0011)
	) read_sdram_0 (
		.clk                  (clk_clk),                                  //         clock.clk
		.reset_n              (~rst_controller_reset_out_reset),          //         reset.reset_n
		.read_en              (read_sdram_read_en),                       //   conduit_end.export
		.data                 (read_sdram_data),                          //              .export
		.addr                 (read_sdram_addr),                          //              .export
		.dev_idle             (read_sdram_dev_idle),                      //              .export
		.data_avalid          (read_sdram_data_avalid),                   //              .export
		.master_waitequest    (read_sdram_0_avalon_master_waitrequest),   // avalon_master.waitrequest
		.master_readdata      (read_sdram_0_avalon_master_readdata),      //              .readdata
		.master_readdatavalid (read_sdram_0_avalon_master_readdatavalid), //              .readdatavalid
		.master_address       (read_sdram_0_avalon_master_address),       //              .address
		.master_byteenable    (read_sdram_0_avalon_master_byteenable),    //              .byteenable
		.master_read          (read_sdram_0_avalon_master_read)           //              .read
	);

	WRITE_SDRAM_FIFO_BURST #(
		.IDLE                 (7'b0000001),
		.START                (7'b0000010),
		.PREPARE_DAT_AND_ADDR (7'b0000100),
		.WRITE_EN             (7'b0001000),
		.WAIT_WRITE_SUCCESS   (7'b0010000),
		.WRITE_SUCCESS        (7'b0100000),
		.BURST_CNT            (6'b010000)
	) write_sdram_burst_0 (
		.clk               (clk_clk),                                       //         clock.clk
		.reset_n           (~rst_controller_reset_out_reset),               //         reset.reset_n
		.write_en          (write_sdram_0_write_en),                        //   conduit_end.export
		.data              (write_sdram_0_data),                            //              .export
		.addr              (write_sdram_0_addr),                            //              .export
		.dev_idle          (write_sdram_0_dev_idle),                        //              .export
		.master_waitequest (write_sdram_burst_0_avalon_master_waitrequest), // avalon_master.waitrequest
		.master_address    (write_sdram_burst_0_avalon_master_address),     //              .address
		.master_byteenable (write_sdram_burst_0_avalon_master_byteenable),  //              .byteenable
		.master_write      (write_sdram_burst_0_avalon_master_write),       //              .write
		.master_writedata  (write_sdram_burst_0_avalon_master_writedata),   //              .writedata
		.master_burstcount (write_sdram_burst_0_avalon_master_burstcount)   //              .burstcount
	);

	WRITE_SDRAM_FIFO_BURST #(
		.IDLE                 (7'b0000001),
		.START                (7'b0000010),
		.PREPARE_DAT_AND_ADDR (7'b0000100),
		.WRITE_EN             (7'b0001000),
		.WAIT_WRITE_SUCCESS   (7'b0010000),
		.WRITE_SUCCESS        (7'b0100000),
		.BURST_CNT            (6'b010000)
	) write_sdram_burst_1 (
		.clk               (clk_clk),                                       //         clock.clk
		.reset_n           (~rst_controller_reset_out_reset),               //         reset.reset_n
		.write_en          (write_sdram_2_1_write_en),                      //   conduit_end.export
		.data              (write_sdram_2_1_data),                          //              .export
		.addr              (write_sdram_2_1_addr),                          //              .export
		.dev_idle          (write_sdram_2_1_dev_idle),                      //              .export
		.master_waitequest (write_sdram_burst_1_avalon_master_waitrequest), // avalon_master.waitrequest
		.master_address    (write_sdram_burst_1_avalon_master_address),     //              .address
		.master_byteenable (write_sdram_burst_1_avalon_master_byteenable),  //              .byteenable
		.master_write      (write_sdram_burst_1_avalon_master_write),       //              .write
		.master_writedata  (write_sdram_burst_1_avalon_master_writedata),   //              .writedata
		.master_burstcount (write_sdram_burst_1_avalon_master_burstcount)   //              .burstcount
	);

	WRITE_SDRAM_FIFO_BURST #(
		.IDLE                 (7'b0000001),
		.START                (7'b0000010),
		.PREPARE_DAT_AND_ADDR (7'b0000100),
		.WRITE_EN             (7'b0001000),
		.WAIT_WRITE_SUCCESS   (7'b0010000),
		.WRITE_SUCCESS        (7'b0100000),
		.BURST_CNT            (6'b010000)
	) write_sdram_burst_2 (
		.clk               (clk_clk),                                       //         clock.clk
		.reset_n           (~rst_controller_reset_out_reset),               //         reset.reset_n
		.write_en          (write_sdram_2_write_en),                        //   conduit_end.export
		.data              (write_sdram_2_data),                            //              .export
		.addr              (write_sdram_2_addr),                            //              .export
		.dev_idle          (write_sdram_2_dev_idle),                        //              .export
		.master_waitequest (write_sdram_burst_2_avalon_master_waitrequest), // avalon_master.waitrequest
		.master_address    (write_sdram_burst_2_avalon_master_address),     //              .address
		.master_byteenable (write_sdram_burst_2_avalon_master_byteenable),  //              .byteenable
		.master_write      (write_sdram_burst_2_avalon_master_write),       //              .write
		.master_writedata  (write_sdram_burst_2_avalon_master_writedata),   //              .writedata
		.master_burstcount (write_sdram_burst_2_avalon_master_burstcount)   //              .burstcount
	);

	sdram_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                       //                                clk_0_clk.clk
		.read_sdram_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // read_sdram_0_reset_reset_bridge_in_reset.reset
		.read_sdram_0_avalon_master_address             (read_sdram_0_avalon_master_address),            //               read_sdram_0_avalon_master.address
		.read_sdram_0_avalon_master_waitrequest         (read_sdram_0_avalon_master_waitrequest),        //                                         .waitrequest
		.read_sdram_0_avalon_master_byteenable          (read_sdram_0_avalon_master_byteenable),         //                                         .byteenable
		.read_sdram_0_avalon_master_read                (read_sdram_0_avalon_master_read),               //                                         .read
		.read_sdram_0_avalon_master_readdata            (read_sdram_0_avalon_master_readdata),           //                                         .readdata
		.read_sdram_0_avalon_master_readdatavalid       (read_sdram_0_avalon_master_readdatavalid),      //                                         .readdatavalid
		.write_sdram_burst_0_avalon_master_address      (write_sdram_burst_0_avalon_master_address),     //        write_sdram_burst_0_avalon_master.address
		.write_sdram_burst_0_avalon_master_waitrequest  (write_sdram_burst_0_avalon_master_waitrequest), //                                         .waitrequest
		.write_sdram_burst_0_avalon_master_burstcount   (write_sdram_burst_0_avalon_master_burstcount),  //                                         .burstcount
		.write_sdram_burst_0_avalon_master_byteenable   (write_sdram_burst_0_avalon_master_byteenable),  //                                         .byteenable
		.write_sdram_burst_0_avalon_master_write        (write_sdram_burst_0_avalon_master_write),       //                                         .write
		.write_sdram_burst_0_avalon_master_writedata    (write_sdram_burst_0_avalon_master_writedata),   //                                         .writedata
		.write_sdram_burst_1_avalon_master_address      (write_sdram_burst_1_avalon_master_address),     //        write_sdram_burst_1_avalon_master.address
		.write_sdram_burst_1_avalon_master_waitrequest  (write_sdram_burst_1_avalon_master_waitrequest), //                                         .waitrequest
		.write_sdram_burst_1_avalon_master_burstcount   (write_sdram_burst_1_avalon_master_burstcount),  //                                         .burstcount
		.write_sdram_burst_1_avalon_master_byteenable   (write_sdram_burst_1_avalon_master_byteenable),  //                                         .byteenable
		.write_sdram_burst_1_avalon_master_write        (write_sdram_burst_1_avalon_master_write),       //                                         .write
		.write_sdram_burst_1_avalon_master_writedata    (write_sdram_burst_1_avalon_master_writedata),   //                                         .writedata
		.write_sdram_burst_2_avalon_master_address      (write_sdram_burst_2_avalon_master_address),     //        write_sdram_burst_2_avalon_master.address
		.write_sdram_burst_2_avalon_master_waitrequest  (write_sdram_burst_2_avalon_master_waitrequest), //                                         .waitrequest
		.write_sdram_burst_2_avalon_master_burstcount   (write_sdram_burst_2_avalon_master_burstcount),  //                                         .burstcount
		.write_sdram_burst_2_avalon_master_byteenable   (write_sdram_burst_2_avalon_master_byteenable),  //                                         .byteenable
		.write_sdram_burst_2_avalon_master_write        (write_sdram_burst_2_avalon_master_write),       //                                         .write
		.write_sdram_burst_2_avalon_master_writedata    (write_sdram_burst_2_avalon_master_writedata),   //                                         .writedata
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),            //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),              //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),               //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),           //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),          //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),         //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),      //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),        //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect)          //                                         .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
