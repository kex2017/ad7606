library verilog;
use verilog.vl_types.all;
entity spi_slave_for_stm32 is
    generic(
        AD_BIT_WIDTH    : integer := 12;
        CHANNEL_NUM     : integer := 3;
        READ_DAT        : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        READ_REG        : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        WRITE_REG       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        IDLE            : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        RW_BIT_DAT      : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        RW_SUCCESS      : vl_logic_vector(0 to 5) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        AD9238_CHA0     : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        AD9238_CHA1     : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        AD9238_CHA2     : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0)
    );
    port(
        clk_100m        : in     vl_logic;
        rst_n           : in     vl_logic;
        ad9238_chip_a_clk: out    vl_logic;
        ad9238_chip_a_dclk: in     vl_logic;
        ad9238_chip_a_data: in     vl_logic_vector;
        ad9238_chip_a_cha1_otr: in     vl_logic;
        ad9238_chip_a_cha2_otr: in     vl_logic;
        ad9238_chip_b_clk: out    vl_logic;
        ad9238_chip_b_dclk: in     vl_logic;
        ad9238_chip_b_data: in     vl_logic_vector;
        ad9238_chip_b_cha1_otr: in     vl_logic;
        ad9238_chip_b_cha2_otr: in     vl_logic;
        spi_sclk_form_stm32: in     vl_logic;
        spi_csn_form_stm32: in     vl_logic;
        spi_mosi_form_stm32: in     vl_logic;
        spi_miso_to_stm32: out    vl_logic;
        sdram_buf0_wdat : out    vl_logic_vector(15 downto 0);
        sdram_buf0_waddr: out    vl_logic_vector(31 downto 0);
        sdram_buf0_wr   : out    vl_logic;
        sdram_buf0_idle : in     vl_logic;
        sdram_buf1_wdat : out    vl_logic_vector(15 downto 0);
        sdram_buf1_waddr: out    vl_logic_vector(31 downto 0);
        sdram_buf1_wr   : out    vl_logic;
        sdram_buf1_idle : in     vl_logic;
        sdram_buf2_wdat : out    vl_logic_vector(15 downto 0);
        sdram_buf2_waddr: out    vl_logic_vector(31 downto 0);
        sdram_buf2_wr   : out    vl_logic;
        sdram_buf2_idle : in     vl_logic;
        sdram_buf_rdat  : in     vl_logic_vector(15 downto 0);
        sdram_buf_raddr : out    vl_logic_vector(31 downto 0);
        sdram_buf_rd    : out    vl_logic;
        sdram_buf_data_avalid: in     vl_logic;
        sdram_idle      : in     vl_logic;
        fpga_interrupt  : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AD_BIT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CHANNEL_NUM : constant is 1;
    attribute mti_svvh_generic_type of READ_DAT : constant is 1;
    attribute mti_svvh_generic_type of READ_REG : constant is 1;
    attribute mti_svvh_generic_type of WRITE_REG : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of RW_BIT_DAT : constant is 1;
    attribute mti_svvh_generic_type of RW_SUCCESS : constant is 1;
    attribute mti_svvh_generic_type of AD9238_CHA0 : constant is 1;
    attribute mti_svvh_generic_type of AD9238_CHA1 : constant is 1;
    attribute mti_svvh_generic_type of AD9238_CHA2 : constant is 1;
end spi_slave_for_stm32;
